module nal

pub fn compile(flags []string) {
	println(flags)
}